library verilog;
use verilog.vl_types.all;
entity ParteAri_vlg_vec_tst is
end ParteAri_vlg_vec_tst;
