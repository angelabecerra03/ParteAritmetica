library verilog;
use verilog.vl_types.all;
entity PartAritmetica is
    port(
        a               : out    vl_logic;
        A0              : in     vl_logic;
        S1              : in     vl_logic;
        A2              : in     vl_logic;
        A1              : in     vl_logic;
        A3              : in     vl_logic;
        S0              : in     vl_logic;
        B0              : in     vl_logic;
        B1              : in     vl_logic;
        B2              : in     vl_logic;
        B3              : in     vl_logic;
        b               : out    vl_logic;
        c               : out    vl_logic;
        d               : out    vl_logic;
        e               : out    vl_logic;
        f               : out    vl_logic;
        g               : out    vl_logic;
        Cout            : out    vl_logic
    );
end PartAritmetica;
