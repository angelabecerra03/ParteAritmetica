library verilog;
use verilog.vl_types.all;
entity FUA_vlg_vec_tst is
end FUA_vlg_vec_tst;
