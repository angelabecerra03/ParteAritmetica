library verilog;
use verilog.vl_types.all;
entity PartAritmetica_vlg_vec_tst is
end PartAritmetica_vlg_vec_tst;
